`ifndef registers_rgu
`define registers_rgu

reg [31:0] RGU_GLB;
reg [31:0] RGU_RST_STATUS;
reg [31:0] RGU_TIMER0;
reg [31:0] RGU_TIMER1;
reg [31:0] RGU_SB_SWRST;
reg [31:0] RGU_SYS_SWRST;
reg [31:0] RGU_SRAM_SWRST;
reg [31:0] RGU_DDR_SWRST;
reg [31:0] RGU_USB_SWRST;
reg [31:0] RGU_MMC_SWRST;
reg [31:0] RGU_DMAC_SWRST;
reg [31:0] RGU_QSPI_SWRST;
reg [31:0] RGU_SPI_SWRST;
reg [31:0] RGU_I2C_SWRST;
reg [31:0] RGU_UART_SWRST;
reg [31:0] RGU_GPIO_SWRST;
reg [31:0] RGU_I2S_SWRST;
reg [31:0] RGU_GPU_SWRST;
reg [31:0] RGU_VIDEC_SWRST;
reg [31:0] RGU_VICOD_SWRST;
reg [31:0] RGU_CAMERA_SWRST;
reg [31:0] RGU_DISPLAY_SWRST;
reg [31:0] RGU_LLC_SWRST;
reg [31:0] RGU_CPU_SWRST;
reg [31:0] RGU_PWM_SWRST ;
reg [31:0] RGU_CPU_PWRUP_SWRST;
reg [31:0] RGU_CPU_PWRUP_HEAVY_­SWRST;

wire SB_DMAC_SWRST;
wire SB_QSPI_SWRST;
wire SB_I2C_SWRST[1:0];
wire SB_UART_SWRST;
wire SB_GPIO_SWRST;
wire SB_SRAM_SWRST;

wire SYS_SWRST;
 
wire SRAM_SWRST;
wire DDR_SWRST;
wire USB_SWRST[3:0];
wire MMC_SWRST[3:0];
wire DMAC_SWRST;
wire QSPI_SWRST[1:0];
wire SPI_SWRST[5:0];
wire I2C_SWRST[6:0];
wire UART_SWRST[4:0];
wire GPIO_SWRST[1:0];
wire I2S_SWRST[1:0];
wire GPU_SWRST;
wire VIDEC_SWRST;
wire VICOD_SWRST;
wire CAMERA_SWRST;
wire DISPLAY_SWRST[1:0];
wire PWM_SWRST[2:0];
wire LLC_SWRST;
wire CPU_SWRST[7:0];
wire CPU_PWRUP_SWRST;
wire CPU_PWRUP_HEAVY_SWRST;


assign SB_DMAC_SWRST = RGU_SB_SWRST[0];
assign SB_QSPI_SWRST = RGU_SB_SWRST[1];
assign SB_I2C_SWRST[1:0] = RGU_SB_SWRST[3:2];
assign SB_UART_SWRST = RGU_SB_SWRST[4];
assign SB_GPIO_SWRST = RGU_SB_SWRST[5];
assign SB_SRAM_SWRST = RGU_SB_SWRST[6];
assign SYS_SWRST = RGU_SYS_SWRST[0];
assign SRAM_SWRST = RGU_SRAM_SWRST[0];
assign DDR_SWRST = RGU_DDR_SWRST[0];
assign USB_SWRST[3:0] = RGU_USB_SWRST[3:0];
assign MMC_SWRST[3:0] = RGU_MMC_SWRST[3:0];
assign DMAC_SWRST = RGU_DMAC_SWRST[0];
assign QSPI_SWRST[1:0] = RGU_QSPI_SWRST[1:0];
assign SPI_SWRST[5:0] = RGU_SPI_SWRST[5:0];
assign I2C_SWRST[6:0] = RGU_I2C_SWRST[6:0];
assign UART_SWRST[4:0] = RGU_UART_SWRST[4:0];
assign GPIO_SWRST[1:0] = RGU_GPIO_SWRST[1:0];
assign I2S_SWRST[1:0] = RGU_I2S_SWRST[1:0];
assign GPU_SWRST = RGU_GPU_SWRST[0];
assign VIDEC_SWRST = RGU_VIDEC_SWRST[0];
assign VICOD_SWRST = RGU_VICOD_SWRST[0];
assign CAMERA_SWRST = RGU_CAMERA_SWRST[0];
assign DISPLAY_SWRST[1:0] = RGU_DISPLAY_SWRST[1:0];
assign PWM_SWRST[2:0] = RGU_PWM_SWRST[2:0];
assign LLC_SWRST = RGU_LLC_SWRST[0];
assign CPU_SWRST[7:0] = RGU_CPU_SWRST[7:0];
assign CPU_PWRUP_SWRST = RGU_CPU_PWRUP_SWRST[0];
assign CPU_PWRUP_HEAVY_SWRST = RGU_CPU_PWRUP_HEAVY_SWRST[0];

// RGU_SB_SWRST.DMAC_SWRST
// RGU_SB_SWRST.QSPI_SWRST
// RGU_SB_SWRST.I2C_SWRST[1:0]
// RGU_SB_SWRST.UART_SWRST
// RGU_SB_SWRST.GPIO_SWRST
// RGU_SB_SWRST.SRAM_SWRST

// RGU_SYS_SWRST.SYS_SWRST

// RGU_SRAM_SWRST.SRAM_SWRST
// RGU_DDR_SWRST.DDR_SWRST
// RGU_USB_SWRST.USB_SWRST[3:0]
// RGU_MMC_SWRST.MMC_SWRST[3:0]
// RGU_DMAC_SWRST.DMAC_SWRST
// RGU_QSPI_SWRST.QSPI_SWRST[1:0]
// RGU_SPI_SWRST.SPI_SWRST[5:0]
// RGU_I2C_SWRST.I2C_SWRST[6:0]
// RGU_UART_SWRST.UART_SWRST[4:0]
// RGU_GPIO_SWRST.GPIO_SWRST[1:0]
// RGU_I2S_SWRST.I2S_SWRST[1:0]
// RGU_GPU_SWRST.GPU_SWRST
// RGU_VIDEC_SWRST.VIDEC_SWRST
// RGU_VICOD_SWRST.VICOD_SWRST
// RGU_CAMERA_SWRST.CAMERA_SWRST
// RGU_DISPLAY_SWRST.DISPLAY_SWRST[1:0]
// RGU_PWM_SWRST.PWM_SWRST[2:0]
// RGU_LLC_SWRST.LLC_SWRST
// RGU_CPU_SWRST.CPU_SWRST[7:0]
// RGU_CPU_PWRUP_SWRST.CPU_PWRUP_SWRST
// RGU_CPU_PWRUP_HEAVY_SWRST.CPU_PWRUP_HEAVY_SWRST
`define RESET_REGS \
RGU_GLB <= 32'h0 ;\
RGU_TIMER0 <= 32'h400 ;\
RGU_TIMER1 <= 32'h400 ;\
RGU_SB_SWRST <= 32'h0 ;\
RGU_SYS_SWRST <= 32'h1 ;\
RGU_SRAM_SWRST <= 32'h1 ;\
RGU_DDR_SWRST <= 32'h1 ;\
RGU_USB_SWRST <= 32'hf ;\
RGU_MMC_SWRST <= 32'hf ;\
RGU_DMAC_SWRST <= 32'h1 ;\
RGU_QSPI_SWRST <= 32'h3 ;\
RGU_SPI_SWRST <= 32'h3f ;\
RGU_I2C_SWRST <= 32'h7f ;\
RGU_UART_SWRST <= 32'h1f ;\
RGU_GPIO_SWRST <= 32'h3 ;\
RGU_I2S_SWRST <= 32'h3 ;\
RGU_GPU_SWRST <= 32'h1 ;\
RGU_VIDEC_SWRST <= 32'h1 ;\
RGU_VICOD_SWRST <= 32'h1;\
RGU_CAMERA_SWRST <= 32'h1 ;\
RGU_DISPLAY_SWRST <= 32'h3 ;\
RGU_LLC_SWRST <= 32'h1 ;\
RGU_CPU_SWRST <= 32'hff ;\
RGU_PWM_SWRST  <= 32'h7f ;\
RGU_CPU_PWRUP_SWRST <= 32'h1 ;\
RGU_CPU_PWRUP_HEAVY_­SWRST <= 32'h1 ;

`endif