module rgu_main(input clk);
    always @(clk) begin
        $display("Hi boss");
    end
endmodule
