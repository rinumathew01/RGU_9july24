interface rgu_intf;
    logic clk;
    logic sys_pwrgd;
    logic sys_reset_n;
    logic sb_wdt_rst_n;
    logic [3:0] wdt_rst_n;
    
    logic rst_sb_sys_n;
    logic rst_sb_dmac_n;
    logic rst_sb_qspi_n;
    logic [1:0] rst_sb_i2c_n;
    logic rst_sb_uart_n;
    logic rst_sb_gpio_n;
    logic rst_sb_sram_n;
    logic rst_sb_wdt_n;
    logic rst_sb_cpu_n;
    logic rst_sys_n;
    logic [3:0] rst_wdt_n;
    logic [7:0] rst_gpt_n;
    logic rst_sram_n;
    logic rst_ddr_n;
    logic [3:0] rst_usb_n;
    logic [3:0] rst_mmc_n;
    logic rst_dmac_n;
    logic [1:0] rst_qspi_n;
    logic [5:0] rst_spi_n;
    logic [6:0] rst_i2c_n;
    logic [4:0] rst_uart_n;
    logic [1:0] rst_gpio_n;
    logic [2:0] rst_pwm_n;
    logic [1:0] rst_i2s_n;
    logic rst_gpu_n;
    logic rst_videc_n;
    logic rst_vicod_n;
    logic [1:0] rst_camera_n;
    logic rst_display_n;
    logic rst_llc_n;
    logic [7:0] rst_cpu_n;
    logic i_test_mode;
    logic i_dft_scan_mode;
    logic i_dft_test_rstn;
endinterface: rgu_intf
