
// Note signal bundle only
interface rgu_if;

  logic clk;
  logic[7:0] cs;
  logic miso;
  logic mosi;
endinterface: rgu_if
