package rgu_test_lib_pkg;

  // Standard UVM import & include:
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  // Any further package imports:
  import rgu_env_pkg::*;
  import apb_agent_pkg::*;
  import rgu_agent_pkg::*;
  import rgu_bus_sequence_lib_pkg::*;
  import rgu_test_seq_lib_pkg::*;
  import rgu_reg_pkg::*;

  // Includes:
`include "rgu_test_base.svh"

endpackage: rgu_test_lib_pkg
